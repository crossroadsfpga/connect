/* =========================================================================
 *
 * Filename:            MCInternalTypes.bsv
 * Date created:        03-16-2011
 * Last modified:       04-06-2011
 * Authors:		Michael Papamichael <papamixATcs.cmu.edu>
 *
 * Description:
 * Types used internally for Memocode network simulator.
 * 
 * =========================================================================
 */

import Vector::*;
import FShow::*;
`include "NetworkExternalTypes.bsv"
//import MCExternalTypes::*;

`include "inc.v"

///////////////////////////////////////////////////////////////////////////////////////////////
// Set network and router parameters
// include *.conf.bsv file generated by running parse_conf on the network configuration file
///////////////////////////////////////////////////////////////////////////////////////////////

//`include "conf_parameters.bsv"
//`include "net_configs/mesh_2x2.txt.conf.bsv"

////////////////////////////////////////////////////////////////////
// Type Definitions
////////////////////////////////////////////////////////////////////
typedef enum{ SepIFRoundRobin, SepOFRoundRobin, SepIFStatic, SepOFStatic, Memocode } AllocType_t deriving(Bits, Eq);

typedef Bit#(n) NumTypeParam#(numeric type n);
// Width of data field in each flit
//typedef 256 FlitDataWidth;
// Max number of flits per packet - check with Derek what the maximum number of flits is - reference uses uchar, i.e. 0-255
typedef 256  MaxNumFlitsPerPacket;
// Max number of traffic entries
typedef 1024 MaxNumTrafficEntries;

typedef 48 MaxCyclesLog;      // Log of maximum number of cycles that can be counted
typedef 48 MaxNumPacketsLog;  // Half of Log of maximum number of packets that each traffic generator can send

// Derived parameters
typedef TSub#(CreditDelay, 1) CreditExtraDelay;

typedef Bit#(TLog#(NumInPorts)) InPort_t;
typedef Bit#(TLog#(NumOutPorts)) OutPort_t;

typedef Bit#(MaxCyclesLog) Cycle_t;
typedef Bit#(MaxNumPacketsLog) NumPackets_t;

typedef struct{
  //Bool            is_head; // turns out this was not needed
  Bool            is_tail; // only required for multi-flit packets
  //RouterID_t      dst;
  UserRecvPortID_t        dst;
  //VC_t            vc; // when flit is sitting in the flitbuffer the VC is implied
  FlitData_t      data; // payload of flit
} FlitBuffer_t
  deriving(Bits, Eq);

typedef struct{
  Flit_t          flit;    // flit
  OutPort_t       out_port; // out_port
} RoutedFlit_t
  deriving(Bits, Eq);


//typedef struct{
//  //Bool            is_head; // turns out this was not needed
//  Bool            is_tail;
//  RouterID_t      dst;
//  VC_t            vc;  
//  FlitData_t      data; // payload of flit
//  `ifdef EN_DBG_REF
//  Bit#(256)        id;  // only used for validation
//  `endif 
//} Flit_t
//  deriving(Bits, Eq);

////////////////////////////////////////////////
// InPort and OutPort interfaces
// Implemented by routers and traffic sources
////////////////////////////////////////////////
//interface InPort;
//  (* always_ready *) method Action putFlit(Maybe#(Flit_t) flit_in);
//  (* always_ready *) method ActionValue#(Credit_t) getCredits;
//endinterface
//
//interface OutPort;
//  (* always_ready *) method ActionValue#(Maybe#(Flit_t)) getFlit();
//  (* always_ready *) method Action putCredits(Credit_t cr_in);
//endinterface
//
//typedef Maybe#(VC_t) Credit_t;  // credits carry VC to which they belong

/////////////////////////////////////////////////
// Traffic Source Types
/////////////////////////////////////////////////
typedef Bit#(TLog#(MaxNumTrafficEntries)) TrafficEntryID_t;
typedef Bit#(TLog#(MaxNumFlitsPerPacket)) FlitID_t;
// Check with Derek what the maximum number of flits is - It is a uchar, i.e. 255
typedef struct{
  RouterID_t        dst;
  VC_t              vc;
  FlitID_t          num_flits;
} TrafficEntry_t
  deriving(Bits, Eq);


//////////////////////////////////////////////////
// Command interface used by MicroBlaze
//////////////////////////////////////////////////

// All possible commands that can be issued through MicroBlaze. 
// Notes: Top module will need to maintain a counter that holds the current TrafficEntryID. This counter 
// needs to get reset using the SetTrafficEntryCount command when starting to populate a new routers traffic entries.

// Used to split cycle values in two halves when bringing in the results through Microblaze 32-bit interface
typedef TDiv#(MaxCyclesLog,2)      HalfMaxCyclesLog;      // Log of maximum number of cycles that can be counted
typedef TDiv#(MaxNumPacketsLog, 2) HalfMaxNumPacketsLog;  // Half of Log of maximum number of packets that each traffic generator can send
typedef Bit#(HalfMaxCyclesLog)     HalfCycle_t;
typedef Bit#(HalfMaxNumPacketsLog) HalfNumPackets_t;

// Command to set current RouterID that will be configured
typedef struct{
  Bit#(8)    rt_id;   // Router ID. Will be truncated to match RouterID_t.
} SetRouterIDCmd_t
  deriving (Bits, Eq);

// Command for setting Route Table entries for currently selected router.
typedef struct{ 
  Bool       endOfTable;  // indicates that route table that was populated should now be committed to BRAM.
  Bit#(8)    dst;         // Destination. Will be truncated to match RouterID_t.
  Bit#(4)    out_p;       // Out Port. Will be truncated to match OutPort_t.
} RouteCmd_t 
  deriving (Bits, Eq);

// Command for setting Traffic Source entries for currently selected router.
typedef struct{ 
  Bool       endOfTraffic;  // indicates end of traffic table for this source. You can commit to BRAM.
  Bit#(8)    dst;        // Destination. Will be truncated to match RouterID_t.
  Bit#(3)    vc;         // VC. Will be truncated to match VC_t.
  Bit#(10)   num_flits;  // Number of flits in packet. Will be truncated to match FlitID_t. 
} TrafficCmd_t
  deriving (Bits, Eq);

// Command for setting Maximum number of packets to be sent by the traffic source of the currently selected router.
// Since MicroBlaze goes through a narrow interface this requires two commands to separately set the high and low halves.
typedef struct{
  Bool              is_lo;           // indicates if this is the lower half of the value.
  HalfNumPackets_t  num_pcks_lo_hi;  // carries low or high half of value.
} SetMaxPcksCmd_t
  deriving (Bits, Eq);

// Command for setting Maximum number of simulation cycles.
// Since MicroBlaze goes through a narrow interface this requires two commands to separately set the high and low halves.
typedef struct{
  Bool              is_lo;
  HalfCycle_t       cycles_lo_hi;
} SetMaxCyclesCmd_t
  deriving (Bits, Eq);

// Command for setting the current traffic entry ID. Only used to set the traffic entry ID to 0, 
// when starting to populate the traffic entries of a new router.
typedef struct{
  TrafficEntryID_t   traf_id;   // Value to set traffic entry ID to. 
} SetTrafficIDCmd_t 
  deriving (Bits, Eq);

// Command wrapper that can contain any of the above commands. This is what the MicroBlaze writes.
typedef union tagged{
    SetRouterIDCmd_t  SetRtID_cmd;
    RouteCmd_t        Route_cmd;
    TrafficCmd_t      Traffic_cmd;
    SetMaxPcksCmd_t   MaxPcks_cmd;
    SetMaxCyclesCmd_t MaxCycles_cmd;
    SetTrafficIDCmd_t SetTrafID_cmd;
    void              InitDone_cmd;
} SetupCmd_t
  deriving (Bits, Eq);

// Results container. Used by MicroBlaze to read simulation results. 
// Since MicroBlaze reads through a narrow interface two commands are require to separately read the high and low halves.
typedef struct{
  Bool           reached_max_cycles;     // indicates if experiment finished because maxCycles where reached
  Bool           is_lo;                  // indicates if this is the lower half of the value.
  HalfCycle_t    elapsed_cycles_lo_hi;   // carries low or high half of value.
} Result_t
  deriving (Bits, Eq);



///////////////////////////////////////////////////
// Data Structures for Virtual Router
///////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////////////////////////////////
// Router state. Includes all state that a router stores and keeps track of, except for route tables.
// Route tables are handled separately, because they have to be initialized by MicroBlaze.
// Used to implement virtual router.
typedef struct{
  //Vector#(NumRouters, OutPort_t)                                        routeTable;
  Vector#(NumInPorts, Vector#(NumVCs, FlitBuffer_t))                    flitBuffers;
  Vector#(NumOutPorts, Vector#(NumVCs, Bool))                           credits;
  Vector#(NumVCs, Vector#(NumInPorts, Vector#(NumOutPorts, Bool)))      hasFlitsVIO;
  Vector#(NumOutPorts, Vector#(NumVCs, Bool ))                          lockedVL;
  Vector#(NumOutPorts, Vector#(NumVCs, InPort_t))                       inPortVL;
} RouterState_t
  deriving (Bits, Eq);

////////////////////////////////////////////////////////////////////////////////////
// Incoming link state. Corresponds to flits and credits going into a router.
typedef struct{
  Vector#(NumInPorts, Maybe#(Flit_t))      in_flits;
  Vector#(NumOutPorts, Credit_t)           in_credits;
} RouterInLinks_t 
  deriving (Bits, Eq);

////////////////////////////////////////////////////////////////////////////////////
// Outgoing link state. Corresponds to flits and credits coming out of a router.
typedef struct{
  Vector#(NumOutPorts, Maybe#(Flit_t))     out_flits;
  Vector#(NumInPorts, Credit_t)            out_credits;
} RouterOutLinks_t
  deriving (Bits, Eq);

///////////////////////////////////////////////////////////////////////////////////////////////////////
// Traffic source state. Includes all state that a traffic source stores and keeps track of.
// Used to implemente virtual traffic source.
typedef struct{
  //Vector#(NumRouters, OutPort_t)                                        routeTable;
  NumPackets_t                     packetsToSend;       // total number of packets to send
  TrafficEntryID_t                 lastTrafficEntryID;  // to know when to wrap-around
  NumPackets_t                     numSentPackets;      // keep track of how many packets have been sent
  TrafficEntry_t                   curTrafficEntry;     // holds current traffic entry
  //TrafficEntryID_t                 curTEindex;          // current Traffic Entry index.
  //FlitID_t                         cur_flits;           // number of flits sent from this packet.
  Vector#(NumVCs, Bool )           credits;             // stores source credits
  // Note: If I uncomment the (wrong) line below the compiler crashes with an internal error message. Send this to Bluespec so they can fix it.
  //Vector#(NumVCs, Reg#(Bool) )     credits;           
} TrafficSourceState_t
  deriving (Bits, Eq);


typedef Bit#(TAdd#( TLog#(NumRouters), TLog#(MaxNumTrafficEntries) ) ) VirtualTrafficEntryID_t;
//typedef Bit#(TLog#(TMul#(NumRouters, MaxNumTrafficEntries))) VirtualTrafficEntryID_t;
//typedef struct{
//  RouterID_t        src_id;    // Traffic Source ID  (one per router)
//  TrafficEntryID_t  traf_id;   // Traffic Entry ID for the traffic table of the specified source
//}  VirtualTrafficEntryID_t
//  deriving (Bits, Eq, Bounded);

interface Network;
  interface Vector#(NumUserSendPorts, InPort)     send_ports;
  interface Vector#(NumUserRecvPorts, OutPort)    recv_ports;
  interface Vector#(NumUserRecvPorts, RecvPortInfo)  recv_ports_info; // Used by clients for obtaining response address
  //interface Vector#(NumRouters, RouterInfo) router_info;
endinterface


///////////////////////////////////////////////////////////////////////////
// Router Interface
interface Router;
  // Port Interfaces
  interface Vector#(NumInPorts, InPort) in_ports;
  interface Vector#(NumOutPorts, OutPort) out_ports;
  // Used to query router info (e.g. ID)
  //interface RouterInfo rt_info;
  //method Action setRoutingEntry(RouterID_t dst, OutPort_t out_p);
endinterface

///////////////////////////////////////////////////////////////////////////
// RouterCore Interface
interface RouterCore;
  interface Vector#(NumInPorts, RouterCoreInPort) in_ports;  // Same as router in_ports, but also carry routing info
  interface Vector#(NumOutPorts, OutPort) out_ports;
  //interface Vector#(NumInPorts, Client#(RouterID_t, OutPort_t)) rt;
endinterface

// InPort interface for RouterCore
interface RouterCoreInPort;
  (* always_ready *) method Action putRoutedFlit(Maybe#(RoutedFlit_t) flit_in);
  (* always_ready *) method ActionValue#(Credit_t) getCredits;
endinterface



interface NetworkSimple;
  interface Vector#(NumUserSendPorts, InPortSimple)     send_ports;
  interface Vector#(NumUserRecvPorts, OutPortSimple)    recv_ports;
  interface Vector#(NumUserRecvPorts, RecvPortInfo)  recv_ports_info; // Used by clients for obtaining response address
  //interface Vector#(NumRouters, RouterInfo) router_info;
endinterface


///////////////////////////////////////////////////////////////////////////
// Router Interface
interface RouterSimple;
  // Port Interfaces
  interface Vector#(NumInPorts, InPortSimple) in_ports;
  interface Vector#(NumOutPorts, OutPortSimple) out_ports;
  // Used to query router info (e.g. ID)
  //interface RouterInfo rt_info;
  //method Action setRoutingEntry(RouterID_t dst, OutPort_t out_p);
endinterface

///////////////////////////////////////////////////////////////////////////
// RouterCore Interface
interface RouterCoreSimple;
  interface Vector#(NumInPorts, RouterCoreInPortSimple) in_ports;  // Same as router in_ports, but also carry routing info
  interface Vector#(NumOutPorts, OutPortSimple) out_ports;
  //interface Vector#(NumInPorts, Client#(RouterID_t, OutPort_t)) rt;
endinterface

// InPort interface for RouterCore
interface RouterCoreInPortSimple;
  (* always_ready *) method Action putRoutedFlit(Maybe#(RoutedFlit_t) flit_in);
  (* always_ready *) method ActionValue#(Vector#(NumVCs, Bool)) getNonFullVCs;
endinterface




/////////////////////////////////////////////////////////////////////////////////
// Add some types to FShow typeclass for pretty printing

instance FShow#(Flit_t);
  function Fmt fshow (Flit_t fl);
    return ($format("Flit [dst:%0d vc:%0d is_tail:%0d data:%x]", fl.dst, fl.vc, fl.is_tail, fl.data));
    //return ($format("Flit [dst:%0d\t vc:%0d\t is_tail:%0d\t data:%x]", fl.dst, fl.vc, fl.is_tail, fl.data));
    //return concatWith("Flit - is_tail:", fshow(""), fshow(fl.is_tail));
    //return concatWith("test"); 
  endfunction
endinstance
