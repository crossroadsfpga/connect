//`define USE_VOQ_ROUTER DEF
`define USE_IQ_ROUTER DEF
`define NUM_USER_SEND_PORTS 16
`define NUM_USER_RECV_PORTS 16
`define NUM_ROUTERS 16
`define NUM_IN_PORTS 5
`define NUM_OUT_PORTS 5
`define CREDIT_DELAY 1
`define NUM_VCS 2
`define ALLOC_TYPE SepIFRoundRobin
`define USE_VIRTUAL_LINKS False
`define FLIT_BUFFER_DEPTH 8
`define FLIT_DATA_WIDTH 32
`define NUM_LINKS 48
`define NETWORK_CUT 0
`define XBAR_LANES 1
`define PIPELINE_CORE False
`define PIPELINE_ALLOCATOR False
`define PIPELINE_LINKS False
